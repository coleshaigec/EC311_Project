module binary_to_BCD(
    input [31:0] thirtytwo_bit_number,
    output [31:0] BCD_number
);
    


endmodule